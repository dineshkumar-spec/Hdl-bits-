module top_module ( input a, input b, output out );
    mod_a inst0(a,b,out);
endmodule
